// draw all triangles on the screen
// draw_start   : trigger signal of drawing
// triangle_data: packed triangle data (projected vertexes on the screen space)
//                [2:0] --- 3 vertexes
//                [1:0] --- x, y coordinates in screen space
//                [9:0] --- 10 bits for each coordinates
// fifo_empty:    indicate whether triangle fifo is empty (so that all triangles are drawn), high when empty
// fifo_r:        read enable signal of triangle fifo, high when read
// DrawX, DrawY:  coordinates of pixels in screen space
// draw_done:     indicate whether drawing is done, high when done
module draw(input Clk, Reset,
            input draw_start,
            input [2:0][1:0][9:0] triangle_data,
            input fifo_empty,
			input [4:0][2:0][35:0] all_proj_vertex,
			input [5:0][5:0] para_out,
			//input [5:0] out1,
            output logic fifo_r,
            output logic [9:0] DrawX, DrawY,
			output logic [23:0]draw_color,
            output logic draw_done
);

    logic draw_triangle_start, draw_triangle_done, draw_surface_start, draw_surface_done;
    logic [1:0][9:0] V1, V2, V3, new_V1, new_V2, new_V3;
	
	logic [9:0] DrawX_T, DrawY_T;
	logic [9:0] DrawX_S, DrawY_S;
	logic [23:0]surface_color;

    // 5 states
    // Wait: wait to start drawing
    // Take1,2: take next triangle data from fifo. 1 for triggering, 2 for taking
    // Draw: draw triangle
    // Done: done	
    enum logic [2:0] {Wait, Take1, Take2, Draw, Surface, Done} curr_state, next_state;
	assign DrawX 		= (curr_state == Surface)?DrawX_S		:DrawX_T;
	assign DrawY 		= (curr_state == Surface)?DrawY_S		:DrawY_T;
	assign draw_color 	= (curr_state == Surface)?surface_color	:{24{(1'b1)}};
	//logic[5:0] para_out;
	//assign para_out=6'b001000;
    // module to draw a triangle
    draw_triangle dl(
                        .Clk(Clk),
                        .Reset(Reset),
                        .draw_triangle_start(draw_triangle_start),
                        .V1(V1),
                        .V2(V2),
                        .V3(V3),
					
                        .DrawX(DrawX_T),
                        .DrawY(DrawY_T),
                        .draw_triangle_done(draw_triangle_done)
						
    );
	point_in ds(
						.Clk(Clk),
                        .Reset(Reset),
						.all_proj_vertex_in(all_proj_vertex),
						.draw_surface_start(draw_surface_start),
						.para_out(para_out),
						.x(DrawX_S),
						.y(DrawY_S),
						.color_out(surface_color),
						.draw_surface_done(draw_surface_done)
	);

    always_ff @(posedge Clk)
    begin
        if (Reset)
        begin
            curr_state <= Done;
            V1 <= 0;
            V2 <= 0;
            V3 <= 0;
        end
        else
        begin
            curr_state <= next_state;
            V1 <= new_V1;
            V2 <= new_V2;
            V3 <= new_V3;
        end
    end

    always_comb
    begin
        next_state = curr_state;
        draw_triangle_start = 1'b0;
		draw_surface_start = 1'b0;
        draw_done = 1'b0;
        fifo_r = 1'b0;
        new_V1 = V1;
        new_V2 = V2;
        new_V3 = V3;
        
        unique case (curr_state)
        Wait:
        begin
            if(draw_start)
                next_state = Take1;
        end
        Take1:
        begin
            if(fifo_empty)
                next_state = Surface;
            else
                next_state = Take2;
        end
        Take2:
        begin
            next_state = Draw;
        end
        Draw:
        begin
            if(draw_triangle_done)
                next_state = Take1;
        end
		Surface:
		begin
			if(draw_surface_done)
				next_state = Done;
		end
        Done:
        begin
            next_state = Wait;
        end
        endcase

        case (curr_state)
        Wait:
        begin
        end
        Take1:
        begin
            fifo_r = 1'b1;
            new_V1 = triangle_data[0];
            new_V2 = triangle_data[1];
            new_V3 = triangle_data[2];
        end
        Take2:
        begin
            new_V1 = triangle_data[0];
            new_V2 = triangle_data[1];
            new_V3 = triangle_data[2];
        end
        Draw:
        begin
            draw_triangle_start = 1'b1;
        end
		Surface:
		begin
			draw_surface_start = 1'b1;
		end
        Done:
        begin
            draw_done = 1'b1;
        end
        endcase
    end

endmodule